// Official code for the Bomberman game, created by Michael Rossinski and Rostyslav Kulnevsky
// 
//
//

module bomberman();

endmodule
	
